module main

import time
import math
import tauraamui.bobatea as tea

struct GameModel {
mut:
	app_send ?fn (tea.Msg)
	window_width int
	window_height int
	position Point
	delta_z  f64 = 1
	frame_label f64
	frame_count int
	last_fps_update time.Time = time.now()
	angle f64
}

struct FrameTickMsg {
	time time.Time
}

fn (mut m GameModel) init() ?tea.Cmd {
	return tea.emit_resize
}

fn (mut m GameModel) update(msg tea.Msg) (tea.Model, ?tea.Cmd) {
	match msg {
		tea.KeyMsg {
			match msg.k_type {
				.special {
					if msg.string() == 'escape' {
						return m.clone(), tea.quit
					}
					match msg.string() {
						'escape' {
							return m.clone(), tea.quit
						}
						else {}
					}
				}
				.runes {
					if msg.string() == 'q' {
						return m.clone(), tea.quit
					}
					if msg.string() == 'x' {
						m.position = Point{ x: m.position.x + 1, y: m.position.y }
						return m.clone(), none
					}
				}
			}
		}
		tea.ResizedMsg {
			m.window_width = msg.window_width
			m.window_height = msg.window_height
		}
		else {}
	}
	return m.clone(), none
}

const vs := [
	Point{x: -0.086914, y: 0.277547, z: 0.400041},
    Point{x: -0.069555, y: 0.329698, z: 0.376422},
    Point{x: -0.125429, y: 0.305056, z: 0.175577},
    Point{x: -0.087431, y: 0.359323, z: 0.182228},
    Point{x: 0.086914, y: 0.277547, z: 0.400041},
    Point{x: 0.069555, y: 0.329698, z: 0.376422},
    Point{x: 0.125429, y: 0.305056, z: 0.175577},
    Point{x: 0.087431, y: 0.359323, z: 0.182228},
    Point{x: -0.162461, y: 0.331177, z: 0.163170},
    Point{x: -0.120032, y: 0.285356, z: 0.287080},
    Point{x: 0.000000, y: 0.316913, z: 0.150254},
    Point{x: 0.000000, y: 0.431152, z: 0.159026},
    Point{x: 0.162461, y: 0.331177, z: 0.163170},
    Point{x: 0.120032, y: 0.285356, z: 0.287080},
    Point{x: 0.038632, y: 0.351515, z: 0.295188},
    Point{x: 0.112575, y: 0.300152, z: 0.416327},
    Point{x: 0.000000, y: 0.283376, z: 0.423906},
    Point{x: 0.000000, y: 0.339429, z: 0.443461},
    Point{x: -0.038632, y: 0.351515, z: 0.295188},
    Point{x: 0.000000, y: 0.333645, z: 0.122512},
    Point{x: 0.151316, y: 0.313187, z: 0.289445},
    Point{x: 0.000000, y: 0.307518, z: 0.456379},
    Point{x: 0.000000, y: 0.299713, z: 0.285755},
    Point{x: 0.000000, y: 0.363275, z: 0.294437},
    Point{x: -0.112575, y: 0.300152, z: 0.416327},
    Point{x: -0.151316, y: 0.313187, z: 0.289445},
    Point{x: 0.118885, y: 0.399961, z: 0.192279},
    Point{x: 0.100036, y: 0.433856, z: 0.198983},
    Point{x: 0.102966, y: 0.396398, z: 0.165539},
    Point{x: 0.084118, y: 0.430293, z: 0.172243},
    Point{x: 0.176608, y: 0.439909, z: 0.152593},
    Point{x: 0.157760, y: 0.473804, z: 0.159297},
    Point{x: 0.160690, y: 0.436346, z: 0.125853},
    Point{x: 0.141841, y: 0.470241, z: 0.132557},
    Point{x: 0.106666, y: 0.390088, z: 0.182523},
    Point{x: 0.104880, y: 0.412922, z: 0.202910},
    Point{x: 0.083687, y: 0.431411, z: 0.190696},
    Point{x: 0.085473, y: 0.408578, z: 0.170310},
    Point{x: 0.132149, y: 0.412268, z: 0.142032},
    Point{x: 0.109170, y: 0.453590, z: 0.150205},
    Point{x: 0.155846, y: 0.457280, z: 0.121927},
    Point{x: 0.177039, y: 0.438791, z: 0.134140},
    Point{x: 0.154060, y: 0.480114, z: 0.142313},
    Point{x: 0.175253, y: 0.461624, z: 0.154527},
    Point{x: 0.151556, y: 0.416612, z: 0.174632},
    Point{x: 0.128577, y: 0.457934, z: 0.182805},
    Point{x: 0.081904, y: 0.401564, z: 0.195735},
    Point{x: 0.116999, y: 0.432110, z: 0.139970},
    Point{x: 0.178822, y: 0.468638, z: 0.129101},
    Point{x: 0.143727, y: 0.438092, z: 0.184867},
    Point{x: 0.146186, y: 0.406646, z: 0.156790},
    Point{x: 0.114539, y: 0.463556, z: 0.168046},
    Point{x: -0.118885, y: 0.399961, z: 0.192279},
    Point{x: -0.100036, y: 0.433856, z: 0.198983},
    Point{x: -0.102966, y: 0.396398, z: 0.165539},
    Point{x: -0.084118, y: 0.430293, z: 0.172243},
    Point{x: -0.176608, y: 0.439909, z: 0.152593},
    Point{x: -0.157760, y: 0.473804, z: 0.159297},
    Point{x: -0.160690, y: 0.436346, z: 0.125853},
    Point{x: -0.141841, y: 0.470241, z: 0.132557},
    Point{x: -0.106666, y: 0.390088, z: 0.182523},
    Point{x: -0.104880, y: 0.412922, z: 0.202910},
    Point{x: -0.083687, y: 0.431411, z: 0.190696},
    Point{x: -0.085473, y: 0.408578, z: 0.170310},
    Point{x: -0.132149, y: 0.412268, z: 0.142032},
    Point{x: -0.109170, y: 0.453590, z: 0.150205},
    Point{x: -0.155846, y: 0.457280, z: 0.121927},
    Point{x: -0.177039, y: 0.438791, z: 0.134140},
    Point{x: -0.154060, y: 0.480114, z: 0.142313},
    Point{x: -0.175253, y: 0.461624, z: 0.154527},
    Point{x: -0.151556, y: 0.416612, z: 0.174632},
    Point{x: -0.128577, y: 0.457934, z: 0.182805},
    Point{x: -0.081904, y: 0.401564, z: 0.195735},
    Point{x: -0.116999, y: 0.432110, z: 0.139970},
    Point{x: -0.178822, y: 0.468638, z: 0.129102},
    Point{x: -0.143727, y: 0.438092, z: 0.184867},
    Point{x: -0.146187, y: 0.406646, z: 0.156790},
    Point{x: -0.114539, y: 0.463556, z: 0.168046},
    Point{x: 0.116485, y: 0.600505, z: 0.141727},
    Point{x: 0.261417, y: -0.299902, z: 0.348366},
    Point{x: -0.116485, y: 0.600505, z: 0.141727},
    Point{x: -0.261417, y: -0.299902, z: 0.348366},
    Point{x: 0.112046, y: 0.657167, z: -0.052576},
    Point{x: 0.239249, y: -0.285613, z: -0.195621},
    Point{x: -0.112046, y: 0.657167, z: -0.052576},
    Point{x: -0.239249, y: -0.285613, z: -0.195621},
    Point{x: 0.182365, y: -0.413886, z: -0.130600},
    Point{x: -0.182365, y: -0.413886, z: -0.130600},
    Point{x: 0.185370, y: -0.411127, z: 0.285766},
    Point{x: -0.185370, y: -0.411127, z: 0.285766},
    Point{x: -0.000000, y: -0.280698, z: -0.288600},
    Point{x: 0.000000, y: 0.685597, z: -0.059119},
    Point{x: -0.000000, y: -0.302354, z: 0.418056},
    Point{x: 0.000000, y: -0.426735, z: -0.175525},
    Point{x: -0.000000, y: 0.616801, z: 0.172179},
    Point{x: 0.346767, y: -0.313945, z: 0.082211},
    Point{x: 0.134460, y: 0.652623, z: 0.053817},
    Point{x: 0.226383, y: -0.434593, z: 0.081386},
    Point{x: 0.000000, y: -0.406050, z: 0.064396},
    Point{x: -0.000000, y: 0.702832, z: 0.076074},
    Point{x: 0.148239, y: 0.499868, z: -0.129503},
    Point{x: 0.167399, y: 0.217376, z: -0.179106},
    Point{x: 0.000000, y: 0.510360, z: -0.177507},
    Point{x: 0.000000, y: 0.222228, z: -0.243510},
    Point{x: 0.000000, y: -0.421023, z: 0.303086},
    Point{x: -0.346767, y: -0.313945, z: 0.082211},
    Point{x: -0.134460, y: 0.652623, z: 0.053817},
    Point{x: 0.253877, y: 0.206739, z: -0.012612},
    Point{x: 0.214625, y: 0.479434, z: 0.003080},
    Point{x: 0.158129, y: 0.450290, z: 0.133907},
    Point{x: 0.188613, y: 0.188153, z: 0.148241},
    Point{x: 0.000000, y: 0.444652, z: 0.202967},
    Point{x: -0.000000, y: 0.189861, z: 0.237317},
    Point{x: -0.226383, y: -0.434593, z: 0.081386},
    Point{x: 0.228074, y: -0.059677, z: -0.205451},
    Point{x: 0.000000, y: -0.055601, z: -0.288645},
    Point{x: -0.000000, y: -0.077669, z: 0.380767},
    Point{x: -0.148239, y: 0.499868, z: -0.129503},
    Point{x: -0.167399, y: 0.217376, z: -0.179106},
    Point{x: 0.336477, y: -0.071376, z: 0.037431},
    Point{x: 0.258730, y: -0.081163, z: 0.294948},
    Point{x: -0.253877, y: 0.206739, z: -0.012612},
    Point{x: -0.214625, y: 0.479434, z: 0.003080},
    Point{x: -0.158129, y: 0.450290, z: 0.133907},
    Point{x: -0.188613, y: 0.188153, z: 0.148241},
    Point{x: -0.228074, y: -0.059677, z: -0.205451},
    Point{x: -0.336477, y: -0.071376, z: 0.037431},
    Point{x: -0.258730, y: -0.081163, z: 0.294948},
    Point{x: 0.066239, y: 0.677571, z: -0.057217},
    Point{x: 0.213490, y: -0.368374, z: -0.165516},
    Point{x: 0.128870, y: -0.280276, z: -0.267035},
    Point{x: 0.106735, y: -0.422750, z: -0.160566},
    Point{x: 0.000000, y: -0.373623, z: -0.249661},
    Point{x: 0.314673, y: -0.301707, z: -0.071136},
    Point{x: -0.314673, y: -0.301707, z: -0.071136},
    Point{x: 0.210922, y: -0.428610, z: -0.043983},
    Point{x: 0.000000, y: -0.423055, z: -0.065328},
    Point{x: -0.244201, y: -0.180778, z: -0.207684},
    Point{x: 0.126667, y: 0.663471, z: -0.006633},
    Point{x: -0.195294, y: 0.491192, z: -0.068821},
    Point{x: 0.000000, y: 0.711143, z: 0.010063},
    Point{x: -0.213490, y: -0.368374, z: -0.165516},
    Point{x: 0.071185, y: 0.691313, z: 0.070402},
    Point{x: -0.155241, y: 0.365055, z: -0.158770},
    Point{x: 0.303068, y: -0.396966, z: 0.087021},
    Point{x: -0.132112, y: 0.602600, z: -0.089009},
    Point{x: 0.120944, y: -0.422690, z: 0.070511},
    Point{x: 0.183037, y: 0.581878, z: 0.028539},
    Point{x: 0.132112, y: 0.602600, z: -0.089009},
    Point{x: 0.155241, y: 0.365055, z: -0.158770},
    Point{x: 0.244201, y: -0.180778, z: -0.207684},
    Point{x: 0.000000, y: 0.617590, z: -0.123992},
    Point{x: 0.000000, y: 0.372508, z: -0.215321},
    Point{x: 0.000000, y: -0.174030, z: -0.298421},
    Point{x: 0.103174, y: 0.187991, z: 0.210662},
    Point{x: 0.000000, y: -0.198444, z: 0.419635},
    Point{x: -0.294693, y: 0.065372, z: 0.007647},
    Point{x: -0.129550, y: 0.627979, z: 0.107967},
    Point{x: 0.294693, y: 0.065372, z: 0.007647},
    Point{x: 0.232020, y: 0.349539, z: -0.013046},
    Point{x: 0.000000, y: 0.323920, z: 0.208490},
    Point{x: 0.088589, y: 0.220688, z: -0.227407},
    Point{x: 0.079730, y: 0.507125, z: -0.165927},
    Point{x: -0.232020, y: 0.349539, z: -0.013046},
    Point{x: 0.195294, y: 0.491192, z: -0.068821},
    Point{x: 0.226314, y: 0.213436, z: -0.101955},
    Point{x: 0.170260, y: 0.326295, z: 0.126748},
    Point{x: -0.000000, y: 0.542220, z: 0.194351},
    Point{x: 0.138605, y: 0.545492, z: 0.141718},
    Point{x: -0.210922, y: -0.428610, z: -0.043983},
    Point{x: 0.224239, y: -0.372873, z: 0.324377},
    Point{x: -0.000000, y: -0.381400, z: 0.379001},
    Point{x: 0.107381, y: -0.417734, z: 0.299738},
    Point{x: 0.069123, y: 0.612108, z: 0.162110},
    Point{x: 0.144110, y: -0.299803, z: 0.404857},
    Point{x: 0.273464, y: -0.200231, z: 0.340419},
    Point{x: 0.086530, y: 0.445098, z: 0.182669},
    Point{x: -0.170260, y: 0.326295, z: 0.126748},
    Point{x: 0.000000, y: 0.670466, z: 0.131824},
    Point{x: -0.226314, y: 0.213436, z: -0.101955},
    Point{x: 0.129550, y: 0.627979, z: 0.107967},
    Point{x: -0.126667, y: 0.663471, z: -0.006633},
    Point{x: 0.240899, y: 0.196199, z: 0.072126},
    Point{x: 0.202094, y: 0.463683, z: 0.072293},
    Point{x: -0.224239, y: -0.372873, z: 0.324377},
    Point{x: 0.196495, y: 0.073973, z: -0.194947},
    Point{x: 0.000000, y: 0.077321, z: -0.268617},
    Point{x: -0.000000, y: 0.053716, z: 0.306623},
    Point{x: 0.356649, y: -0.201172, z: 0.064475},
    Point{x: 0.223708, y: 0.050083, z: 0.216822},
    Point{x: 0.302413, y: -0.064867, z: -0.098045},
    Point{x: -0.138605, y: 0.545492, z: 0.141718},
    Point{x: 0.143359, y: -0.079578, z: 0.361124},
    Point{x: -0.273464, y: -0.200231, z: 0.340419},
    Point{x: 0.122283, y: -0.056588, z: -0.268697},
    Point{x: 0.323489, y: -0.077819, z: 0.178606},
    Point{x: -0.183037, y: 0.581878, z: 0.028539},
    Point{x: 0.211567, y: -0.425514, z: 0.204949},
    Point{x: 0.329913, y: -0.309199, z: 0.232998},
    Point{x: -0.303068, y: -0.396966, z: 0.087021},
    Point{x: 0.000000, y: -0.416129, z: 0.193289},
    Point{x: -0.240899, y: 0.196199, z: 0.072126},
    Point{x: -0.202094, y: 0.463683, z: 0.072293},
    Point{x: -0.196495, y: 0.073973, z: -0.194947},
    Point{x: -0.356649, y: -0.201172, z: 0.064475},
    Point{x: -0.223708, y: 0.050083, z: 0.216822},
    Point{x: -0.302413, y: -0.064867, z: -0.098045},
    Point{x: -0.323489, y: -0.077819, z: 0.178606},
    Point{x: -0.211567, y: -0.425514, z: 0.204949},
    Point{x: -0.329913, y: -0.309199, z: 0.232998},
    Point{x: -0.120944, y: -0.422690, z: 0.070511},
    Point{x: -0.128870, y: -0.280276, z: -0.267035},
    Point{x: -0.106735, y: -0.422750, z: -0.160566},
    Point{x: -0.071185, y: 0.691312, z: 0.070402},
    Point{x: -0.103174, y: 0.187991, z: 0.210662},
    Point{x: -0.144110, y: -0.299803, z: 0.404857},
    Point{x: -0.066239, y: 0.677571, z: -0.057217},
    Point{x: -0.079730, y: 0.507125, z: -0.165927},
    Point{x: -0.088589, y: 0.220688, z: -0.227407},
    Point{x: -0.069123, y: 0.612108, z: 0.162110},
    Point{x: -0.107381, y: -0.417734, z: 0.299738},
    Point{x: -0.086530, y: 0.445098, z: 0.182669},
    Point{x: -0.143359, y: -0.079578, z: 0.361124},
    Point{x: -0.122283, y: -0.056588, z: -0.268697},
    Point{x: -0.116187, y: -0.369086, z: -0.229604},
    Point{x: -0.072661, y: 0.612795, z: -0.116367},
    Point{x: 0.116187, y: -0.369087, z: -0.229604},
    Point{x: 0.113112, y: -0.424606, z: 0.196042},
    Point{x: 0.218688, y: 0.336754, z: 0.060131},
    Point{x: -0.082517, y: 0.370222, z: -0.201199},
    Point{x: -0.342146, y: -0.202745, z: 0.218515},
    Point{x: -0.277483, y: -0.384780, z: -0.052960},
    Point{x: 0.342146, y: -0.202745, z: 0.218515},
    Point{x: -0.123321, y: 0.051288, z: 0.282574},
    Point{x: 0.104612, y: 0.076285, z: -0.250504},
    Point{x: -0.263362, y: 0.070961, z: -0.103638},
    Point{x: 0.072661, y: 0.612795, z: -0.116367},
    Point{x: 0.068288, y: 0.700296, z: 0.006932},
    Point{x: -0.218688, y: 0.336754, z: 0.060131},
    Point{x: -0.068288, y: 0.700296, z: 0.006932},
    Point{x: 0.092843, y: 0.323418, z: 0.183578},
    Point{x: 0.277483, y: -0.384780, z: -0.052960},
    Point{x: -0.092843, y: 0.323418, z: 0.183578},
    Point{x: 0.114344, y: -0.430659, z: -0.055794},
    Point{x: -0.069793, y: 0.661151, z: 0.124576},
    Point{x: 0.123321, y: 0.051288, z: 0.282574},
    Point{x: -0.113112, y: -0.424606, z: 0.196042},
    Point{x: 0.123369, y: -0.375786, z: 0.369703},
    Point{x: 0.069793, y: 0.661151, z: 0.124576},
    Point{x: -0.169024, y: 0.594663, z: -0.036361},
    Point{x: -0.151487, y: -0.198724, z: 0.403451},
    Point{x: 0.082517, y: 0.370222, z: -0.201199},
    Point{x: 0.284665, y: -0.386757, z: 0.223581},
    Point{x: -0.284665, y: -0.386757, z: 0.223581},
    Point{x: -0.077124, y: 0.541621, z: 0.179388},
    Point{x: -0.123369, y: -0.375786, z: 0.369703},
    Point{x: 0.322028, y: -0.191732, z: -0.086948},
    Point{x: -0.114344, y: -0.430659, z: -0.055794},
    Point{x: 0.169024, y: 0.594663, z: -0.036361},
    Point{x: 0.208363, y: 0.358708, z: -0.090994},
    Point{x: 0.077124, y: 0.541621, z: 0.179388},
    Point{x: -0.322028, y: -0.191732, z: -0.086948},
    Point{x: 0.173487, y: 0.562450, z: 0.090260},
    Point{x: 0.263362, y: 0.070961, z: -0.103638},
    Point{x: -0.173487, y: 0.562450, z: 0.090260},
    Point{x: -0.131368, y: -0.175217, z: -0.277201},
    Point{x: -0.208363, y: 0.358708, z: -0.090994},
    Point{x: 0.151487, y: -0.198724, z: 0.403451},
    Point{x: -0.282070, y: 0.056411, z: 0.120093},
    Point{x: 0.131368, y: -0.175217, z: -0.277201},
    Point{x: 0.282071, y: 0.056411, z: 0.120093},
    Point{x: -0.104612, y: 0.076285, z: -0.250504},
    Point{x: -0.508828, y: -0.488737, z: 0.156039},
    Point{x: -0.522541, y: -0.410065, z: 0.161508},
    Point{x: -0.282585, y: -0.488737, z: -0.115427},
    Point{x: -0.282585, y: -0.309773, z: -0.115427},
    Point{x: -0.361756, y: -0.488737, z: 0.278610},
    Point{x: -0.364664, y: -0.410065, z: 0.293084},
    Point{x: -0.135514, y: -0.488737, z: 0.007144},
    Point{x: -0.135514, y: -0.309773, z: 0.007144},
    Point{x: -0.411821, y: -0.495733, z: 0.006876},
    Point{x: -0.549731, y: -0.455582, z: 0.172353},
    Point{x: -0.411821, y: -0.288796, z: 0.006876},
    Point{x: -0.273911, y: -0.455582, z: -0.158601},
    Point{x: -0.184261, y: -0.495733, z: -0.083886},
    Point{x: -0.184261, y: -0.288796, z: -0.083886},
    Point{x: -0.094610, y: -0.455582, z: -0.009170},
    Point{x: -0.232520, y: -0.495733, z: 0.156307},
    Point{x: -0.232520, y: -0.288796, z: 0.156307},
    Point{x: -0.370430, y: -0.455582, z: 0.321783},
    Point{x: -0.460081, y: -0.495733, z: 0.247068},
    Point{x: -0.477521, y: -0.396120, z: 0.267995},
    Point{x: -0.445638, y: -0.455582, z: -0.021308},
    Point{x: -0.132239, y: -0.455582, z: -0.146306},
    Point{x: -0.198703, y: -0.455582, z: 0.184490},
    Point{x: -0.512102, y: -0.455582, z: 0.309488},
    Point{x: -0.322171, y: -0.510414, z: 0.081591},
    Point{x: -0.322171, y: -0.244774, z: 0.081591},
    Point{x: 0.508827, y: -0.488737, z: 0.156039},
    Point{x: 0.522541, y: -0.410065, z: 0.161508},
    Point{x: 0.282585, y: -0.488737, z: -0.115427},
    Point{x: 0.282585, y: -0.309773, z: -0.115427},
    Point{x: 0.361756, y: -0.488737, z: 0.278610},
    Point{x: 0.364664, y: -0.410065, z: 0.293084},
    Point{x: 0.135514, y: -0.488737, z: 0.007144},
    Point{x: 0.135514, y: -0.309773, z: 0.007144},
    Point{x: 0.411821, y: -0.495733, z: 0.006876},
    Point{x: 0.549731, y: -0.455582, z: 0.172353},
    Point{x: 0.411821, y: -0.288796, z: 0.006876},
    Point{x: 0.273911, y: -0.455582, z: -0.158601},
    Point{x: 0.184261, y: -0.495733, z: -0.083886},
    Point{x: 0.184261, y: -0.288796, z: -0.083886},
    Point{x: 0.094610, y: -0.455582, z: -0.009170},
    Point{x: 0.232520, y: -0.495733, z: 0.156307},
    Point{x: 0.232520, y: -0.288796, z: 0.156307},
    Point{x: 0.370430, y: -0.455582, z: 0.321783},
    Point{x: 0.460080, y: -0.495733, z: 0.247068},
    Point{x: 0.477521, y: -0.396120, z: 0.267995},
    Point{x: 0.445638, y: -0.455582, z: -0.021308},
    Point{x: 0.132239, y: -0.455582, z: -0.146306},
    Point{x: 0.198703, y: -0.455582, z: 0.184490},
    Point{x: 0.512102, y: -0.455582, z: 0.309488},
    Point{x: 0.322171, y: -0.510414, z: 0.081591},
    Point{x: 0.322171, y: -0.244774, z: 0.081591},

]

const fs := [
	[22, 2, 10],
    [21, 1, 24],
    [7, 23, 14],
    [2, 25, 8],
    [0, 21, 24],
    [1, 23, 18],
    [3, 23, 11],
    [2, 19, 10],
    [19, 7, 12],
    [6, 19, 12],
    [22, 0, 9],
    [20, 5, 15],
    [13, 15, 4],
    [7, 20, 12],
    [5, 23, 17],
    [25, 1, 18],
    [22, 4, 16],
    [6, 22, 10],
    [19, 3, 11],
    [24, 9, 0],
    [4, 21, 16],
    [5, 21, 15],
    [25, 3, 8],
    [6, 20, 13],
    [34, 35, 46],
    [35, 36, 46],
    [33, 51, 42],
    [36, 37, 46],
    [34, 37, 28],
    [76, 58, 64],
    [28, 50, 34],
    [77, 53, 62],
    [47, 33, 40],
    [76, 52, 70],
    [32, 47, 40],
    [75, 52, 61],
    [28, 47, 38],
    [42, 43, 48],
    [41, 43, 30],
    [40, 42, 48],
    [31, 51, 45],
    [73, 54, 64],
    [50, 30, 44],
    [32, 50, 38],
    [76, 56, 67],
    [75, 53, 71],
    [60, 61, 52],
    [73, 55, 63],
    [61, 62, 53],
    [75, 57, 69],
    [62, 63, 55],
    [77, 55, 65],
    [60, 63, 72],
    [76, 54, 60],
    [59, 73, 66],
    [77, 59, 68],
    [73, 58, 66],
    [29, 47, 37],
    [68, 69, 57],
    [77, 57, 71],
    [67, 69, 74],
    [68, 66, 74],
    [27, 49, 45],
    [75, 56, 70],
    [67, 66, 58],
    [26, 50, 44],
    [49, 26, 44],
    [29, 51, 39],
    [30, 49, 44],
    [31, 49, 43],
    [51, 27, 45],
    [40, 41, 32],
    [90, 224, 211],
    [93, 224, 132],
    [212, 141, 224],
    [224, 85, 211],
    [102, 225, 151],
    [217, 145, 225],
    [225, 84, 216],
    [151, 216, 91],
    [90, 226, 132],
    [83, 226, 130],
    [129, 131, 226],
    [226, 93, 132],
    [88, 227, 197],
    [172, 200, 227],
    [200, 146, 227],
    [227, 97, 197],
    [183, 159, 108],
    [109, 228, 183],
    [166, 182, 228],
    [228, 107, 159],
    [103, 229, 152],
    [218, 143, 229],
    [143, 217, 229],
    [152, 217, 102],
    [204, 207, 126],
    [105, 230, 204],
    [209, 193, 230],
    [230, 127, 207],
    [141, 134, 85],
    [87, 231, 141],
    [231, 113, 199],
    [231, 105, 134],
    [195, 188, 119],
    [120, 232, 195],
    [175, 198, 232],
    [232, 95, 188],
    [187, 222, 116],
    [112, 233, 187],
    [214, 205, 233],
    [233, 127, 222],
    [115, 234, 194],
    [186, 161, 234],
    [234, 101, 185],
    [194, 185, 114],
    [121, 235, 156],
    [179, 203, 235],
    [235, 125, 206],
    [156, 206, 126],
    [102, 236, 162],
    [151, 128, 236],
    [236, 82, 148],
    [162, 148, 100],
    [96, 237, 142],
    [138, 128, 237],
    [237, 91, 140],
    [142, 140, 99],
    [163, 202, 122],
    [121, 238, 163],
    [201, 177, 238],
    [238, 123, 202],
    [106, 239, 181],
    [213, 140, 239],
    [239, 91, 216],
    [181, 216, 84],
    [154, 160, 112],
    [110, 240, 154],
    [240, 109, 176],
    [160, 176, 111],
    [133, 129, 83],
    [95, 241, 133],
    [241, 97, 135],
    [241, 86, 129],
    [160, 214, 112],
    [160, 221, 242],
    [242, 123, 177],
    [242, 124, 214],
    [86, 243, 131],
    [135, 146, 243],
    [243, 98, 136],
    [131, 136, 93],
    [157, 213, 106],
    [80, 244, 157],
    [219, 178, 244],
    [244, 99, 213],
    [192, 187, 116],
    [120, 245, 192],
    [189, 154, 245],
    [245, 112, 187],
    [89, 246, 220],
    [113, 246, 208],
    [210, 200, 246],
    [220, 200, 104],
    [92, 247, 174],
    [171, 172, 247],
    [247, 88, 170],
    [174, 170, 79],
    [142, 180, 96],
    [99, 248, 142],
    [178, 173, 248],
    [248, 78, 180],
    [181, 196, 106],
    [84, 249, 181],
    [145, 139, 249],
    [249, 122, 196],
    [155, 215, 92],
    [155, 222, 250],
    [222, 193, 250],
    [250, 81, 215],
    [103, 251, 161],
    [152, 162, 251],
    [162, 149, 251],
    [161, 149, 101],
    [170, 198, 79],
    [88, 252, 170],
    [197, 144, 252],
    [252, 95, 198],
    [209, 184, 81],
    [105, 253, 209],
    [199, 208, 253],
    [253, 89, 184],
    [111, 254, 221],
    [167, 219, 254],
    [254, 80, 191],
    [221, 191, 123],
    [92, 255, 171],
    [215, 184, 255],
    [255, 89, 220],
    [171, 220, 104],
    [119, 256, 190],
    [188, 133, 256],
    [256, 83, 150],
    [190, 150, 114],
    [87, 257, 169],
    [212, 136, 257],
    [257, 98, 210],
    [169, 210, 113],
    [147, 138, 96],
    [108, 258, 147],
    [164, 148, 258],
    [258, 82, 138],
    [108, 259, 164],
    [159, 165, 259],
    [259, 101, 149],
    [259, 100, 164],
    [111, 260, 167],
    [176, 168, 260],
    [260, 78, 173],
    [167, 173, 94],
    [126, 261, 204],
    [206, 137, 261],
    [261, 85, 134],
    [204, 134, 105],
    [96, 262, 147],
    [78, 262, 180],
    [262, 109, 183],
    [262, 108, 147],
    [107, 263, 165],
    [158, 190, 263],
    [263, 114, 185],
    [165, 185, 101],
    [106, 264, 157],
    [122, 264, 196],
    [264, 123, 191],
    [264, 80, 157],
    [90, 265, 153],
    [211, 137, 265],
    [265, 125, 223],
    [153, 223, 115],
    [122, 266, 163],
    [117, 266, 139],
    [266, 118, 179],
    [163, 179, 121],
    [174, 155, 92],
    [79, 267, 174],
    [175, 192, 267],
    [155, 192, 116],
    [156, 201, 121],
    [126, 268, 156],
    [207, 205, 268],
    [268, 124, 201],
    [90, 269, 130],
    [153, 194, 269],
    [269, 114, 150],
    [130, 150, 83],
    [182, 158, 107],
    [110, 270, 182],
    [189, 195, 270],
    [270, 119, 158],
    [115, 271, 186],
    [223, 203, 271],
    [271, 118, 218],
    [186, 218, 103],
    [272, 292, 280],
    [273, 292, 281],
    [292, 275, 283],
    [292, 274, 280],
    [283, 284, 274],
    [283, 285, 293],
    [285, 286, 293],
    [284, 286, 278],
    [278, 294, 287],
    [279, 294, 286],
    [294, 277, 289],
    [294, 276, 287],
    [289, 290, 276],
    [289, 291, 295],
    [291, 281, 295],
    [290, 281, 272],
    [274, 296, 280],
    [278, 296, 284],
    [296, 276, 290],
    [296, 272, 280],
    [279, 297, 288],
    [275, 297, 285],
    [297, 273, 291],
    [297, 277, 288],
    [298, 318, 307],
    [318, 299, 307],
    [318, 301, 308],
    [300, 318, 306],
    [310, 309, 300],
    [309, 311, 301],
    [312, 311, 319],
    [310, 312, 319],
    [304, 320, 312],
    [320, 305, 312],
    [320, 303, 314],
    [302, 320, 313],
    [316, 315, 302],
    [315, 317, 303],
    [307, 317, 321],
    [316, 307, 321],
    [300, 322, 310],
    [322, 304, 310],
    [322, 302, 313],
    [298, 322, 306],
    [305, 323, 311],
    [323, 301, 311],
    [323, 299, 308],
    [303, 323, 314],
    [22, 9, 2],
    [21, 17, 1],
    [7, 11, 23],
    [2, 9, 25],
    [0, 16, 21],
    [1, 17, 23],
    [3, 18, 23],
    [2, 8, 19],
    [19, 11, 7],
    [6, 10, 19],
    [22, 16, 0],
    [20, 14, 5],
    [13, 20, 15],
    [7, 14, 20],
    [5, 14, 23],
    [25, 24, 1],
    [22, 13, 4],
    [6, 13, 22],
    [19, 8, 3],
    [24, 25, 9],
    [4, 15, 21],
    [5, 17, 21],
    [25, 18, 3],
    [6, 12, 20],
    [34, 26, 35],
    [35, 27, 36],
    [33, 39, 51],
    [36, 29, 37],
    [34, 46, 37],
    [76, 67, 58],
    [28, 38, 50],
    [77, 71, 53],
    [47, 39, 33],
    [76, 60, 52],
    [32, 38, 47],
    [75, 70, 52],
    [28, 37, 47],
    [42, 31, 43],
    [41, 48, 43],
    [40, 33, 42],
    [31, 42, 51],
    [73, 63, 54],
    [50, 41, 30],
    [32, 41, 50],
    [76, 70, 56],
    [75, 61, 53],
    [60, 72, 61],
    [73, 65, 55],
    [61, 72, 62],
    [75, 71, 57],
    [62, 72, 63],
    [77, 62, 55],
    [60, 54, 63],
    [76, 64, 54],
    [59, 65, 73],
    [77, 65, 59],
    [73, 64, 58],
    [29, 39, 47],
    [68, 74, 69],
    [77, 68, 57],
    [67, 56, 69],
    [68, 59, 66],
    [27, 35, 49],
    [75, 69, 56],
    [67, 74, 66],
    [26, 34, 50],
    [49, 35, 26],
    [29, 36, 51],
    [30, 43, 49],
    [31, 45, 49],
    [51, 36, 27],
    [40, 48, 41],
    [90, 132, 224],
    [93, 212, 224],
    [212, 87, 141],
    [224, 141, 85],
    [102, 217, 225],
    [217, 117, 145],
    [225, 145, 84],
    [151, 225, 216],
    [90, 130, 226],
    [83, 129, 226],
    [129, 86, 131],
    [226, 131, 93],
    [88, 172, 227],
    [172, 104, 200],
    [200, 98, 146],
    [227, 146, 97],
    [183, 228, 159],
    [109, 166, 228],
    [166, 110, 182],
    [228, 182, 107],
    [103, 218, 229],
    [218, 118, 143],
    [143, 117, 217],
    [152, 229, 217],
    [204, 230, 207],
    [105, 209, 230],
    [209, 81, 193],
    [230, 193, 127],
    [141, 231, 134],
    [87, 169, 231],
    [231, 169, 113],
    [231, 199, 105],
    [195, 232, 188],
    [120, 175, 232],
    [175, 79, 198],
    [232, 198, 95],
    [187, 233, 222],
    [112, 214, 233],
    [214, 124, 205],
    [233, 205, 127],
    [115, 186, 234],
    [186, 103, 161],
    [234, 161, 101],
    [194, 234, 185],
    [121, 179, 235],
    [179, 118, 203],
    [235, 203, 125],
    [156, 235, 206],
    [102, 151, 236],
    [151, 91, 128],
    [236, 128, 82],
    [162, 236, 148],
    [96, 138, 237],
    [138, 82, 128],
    [237, 128, 91],
    [142, 237, 140],
    [163, 238, 202],
    [121, 201, 238],
    [201, 124, 177],
    [238, 177, 123],
    [106, 213, 239],
    [213, 99, 140],
    [239, 140, 91],
    [181, 239, 216],
    [154, 240, 160],
    [110, 166, 240],
    [240, 166, 109],
    [160, 240, 176],
    [133, 241, 129],
    [95, 144, 241],
    [241, 144, 97],
    [241, 135, 86],
    [160, 242, 214],
    [160, 111, 221],
    [242, 221, 123],
    [242, 177, 124],
    [86, 135, 243],
    [135, 97, 146],
    [243, 146, 98],
    [131, 243, 136],
    [157, 244, 213],
    [80, 219, 244],
    [219, 94, 178],
    [244, 178, 99],
    [192, 245, 187],
    [120, 189, 245],
    [189, 110, 154],
    [245, 154, 112],
    [89, 208, 246],
    [113, 210, 246],
    [210, 98, 200],
    [220, 246, 200],
    [92, 171, 247],
    [171, 104, 172],
    [247, 172, 88],
    [174, 247, 170],
    [142, 248, 180],
    [99, 178, 248],
    [178, 94, 173],
    [248, 173, 78],
    [181, 249, 196],
    [84, 145, 249],
    [145, 117, 139],
    [249, 139, 122],
    [155, 250, 215],
    [155, 116, 222],
    [222, 127, 193],
    [250, 193, 81],
    [103, 152, 251],
    [152, 102, 162],
    [162, 100, 149],
    [161, 251, 149],
    [170, 252, 198],
    [88, 197, 252],
    [197, 97, 144],
    [252, 144, 95],
    [209, 253, 184],
    [105, 199, 253],
    [199, 113, 208],
    [253, 208, 89],
    [111, 167, 254],
    [167, 94, 219],
    [254, 219, 80],
    [221, 254, 191],
    [92, 215, 255],
    [215, 81, 184],
    [255, 184, 89],
    [171, 255, 220],
    [119, 188, 256],
    [188, 95, 133],
    [256, 133, 83],
    [190, 256, 150],
    [87, 212, 257],
    [212, 93, 136],
    [257, 136, 98],
    [169, 257, 210],
    [147, 258, 138],
    [108, 164, 258],
    [164, 100, 148],
    [258, 148, 82],
    [108, 159, 259],
    [159, 107, 165],
    [259, 165, 101],
    [259, 149, 100],
    [111, 176, 260],
    [176, 109, 168],
    [260, 168, 78],
    [167, 260, 173],
    [126, 206, 261],
    [206, 125, 137],
    [261, 137, 85],
    [204, 261, 134],
    [96, 180, 262],
    [78, 168, 262],
    [262, 168, 109],
    [262, 183, 108],
    [107, 158, 263],
    [158, 119, 190],
    [263, 190, 114],
    [165, 263, 185],
    [106, 196, 264],
    [122, 202, 264],
    [264, 202, 123],
    [264, 191, 80],
    [90, 211, 265],
    [211, 85, 137],
    [265, 137, 125],
    [153, 265, 223],
    [122, 139, 266],
    [117, 143, 266],
    [266, 143, 118],
    [163, 266, 179],
    [174, 267, 155],
    [79, 175, 267],
    [175, 120, 192],
    [155, 267, 192],
    [156, 268, 201],
    [126, 207, 268],
    [207, 127, 205],
    [268, 205, 124],
    [90, 153, 269],
    [153, 115, 194],
    [269, 194, 114],
    [130, 269, 150],
    [182, 270, 158],
    [110, 189, 270],
    [189, 120, 195],
    [270, 195, 119],
    [115, 223, 271],
    [223, 125, 203],
    [271, 203, 118],
    [186, 271, 218],
    [272, 281, 292],
    [273, 282, 292],
    [292, 282, 275],
    [292, 283, 274],
    [283, 293, 284],
    [283, 275, 285],
    [285, 279, 286],
    [284, 293, 286],
    [278, 286, 294],
    [279, 288, 294],
    [294, 288, 277],
    [294, 289, 276],
    [289, 295, 290],
    [289, 277, 291],
    [291, 273, 281],
    [290, 295, 281],
    [274, 284, 296],
    [278, 287, 296],
    [296, 287, 276],
    [296, 290, 272],
    [279, 285, 297],
    [275, 282, 297],
    [297, 282, 273],
    [297, 291, 277],
    [298, 306, 318],
    [318, 308, 299],
    [318, 309, 301],
    [300, 309, 318],
    [310, 319, 309],
    [309, 319, 311],
    [312, 305, 311],
    [310, 304, 312],
    [304, 313, 320],
    [320, 314, 305],
    [320, 315, 303],
    [302, 315, 320],
    [316, 321, 315],
    [315, 321, 317],
    [307, 299, 317],
    [316, 298, 307],
    [300, 306, 322],
    [322, 313, 304],
    [322, 316, 302],
    [298, 316, 322],
    [305, 314, 323],
    [323, 308, 301],
    [323, 317, 299],
    [303, 317, 323],
]

fn translate_z(p Point, delta_z f64) Point {
	return Point{
		x: p.x
		y: p.y
		z: p.z + delta_z
	}
}

fn rotate_xz(p Point, angle f64) Point {
	c := math.cos(angle)
	s := math.sin(angle)
	return Point{
		x: (p.x * c) - (p.z * s)
		y: p.y
		z: (p.z * s) + (p.z * c)
	}
}

fn (mut m GameModel) view(mut ctx tea.Context) {
	// m.delta_z += (m.frame_label / 1000.0)
	m.angle += math.pi * (m.frame_label / 1000.0)

	ctx.set_bg_color(tea.Color{ 30, 30, 30 })
	ctx.draw_rect(0, 0, m.window_width, m.window_height)
	ctx.reset_bg_color()

	ctx.set_bg_color(tea.Color{ g: 200 })

	/*
	for v in vs {
		point(mut ctx, screen(m.window_width, m.window_height, project(translate_z(rotate_xz(v, m.angle), m.delta_z))))
	}
	*/

	for f in fs {
		for i in 0..f.len {
			a := vs[f[i]]
			b := vs[f[(i + 1) % f.len]]
			line(mut ctx, screen(m.window_width, m.window_height, project(translate_z(rotate_xz(a, m.angle), m.delta_z))),
			screen(m.window_width, m.window_height, project(translate_z(rotate_xz(b, m.angle), m.delta_z))))
		}
	}

	ctx.reset_bg_color()

	ctx.set_color(tea.Color.ansi(255))
	ctx.draw_text(1, 1, "frames: ${m.frame_label}, DELTA Z: ${1 + m.delta_z}")

	if time.now() - m.last_fps_update >= (1 * time.second) {
		m.frame_label = 1000.0 / f64(m.frame_count)
		m.frame_count = 0
		m.last_fps_update = time.now()
	}
	m.frame_count += 1
}

fn (m GameModel) clone() tea.Model {
	return GameModel{
		...m
	}
}

struct Point{
	x f64
	y f64
	z f64
}

fn point(mut ctx tea.Context, p Point) {
	s := 1.0
	ctx.draw_rect(int(p.x - s / 2), int(p.y - s / 2), int(s), int(s))
}

fn line(mut ctx tea.Context, p1 Point, p2 Point) {
	ctx.draw_line(int(p1.x), int(p1.y), int(p2.x), int(p2.y), false)
}

fn screen(width int, height int, p Point) Point {
	w := f64(width)
	h := f64(height)
	return Point{
		x: (p.x + 1) / 2 * w
		y: (1 - (p.y + 1) / 2) * h
	}
}

fn project(p Point) Point {
	return Point{
		x: p.x / p.z
		y: p.y / p.z
	}
}

fn main() {
	mut game_model := GameModel{}
	mut app := tea.new_program(mut game_model)
	game_model.app_send = app.send
	app.run() or { panic('something went wrong! ${err}') }
}

